module top ( 
	) ;

